module top ( 
	) ;

